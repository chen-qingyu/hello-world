// Verilog
// Icarus Verilog version 12.0

module main();
    initial begin
        $display("Hello World!");
    end
endmodule
