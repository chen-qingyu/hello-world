// Verilog
// Icarus Verilog version 12.0
// iverilog -o HelloWorld HelloWorld.v; vvp HelloWorld

module main();
    initial begin
        $display("Hello World!");
    end
endmodule
